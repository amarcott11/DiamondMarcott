module datapath(input)



endmodule